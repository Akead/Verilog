module fun(input [2:0] A, input [2:0] B, output C, D);

	assign C = (~B[1] & ~B[0] & ~A[2] & A[0]) | (~B[1] & ~A[2] & A[1]) | (~B[0] & ~A[2] & A[1] & A[0]) | (B[2] & ~A[2]) | (B[2] & ~B[1] & ~B[0] & A[0]) | (B[2] & ~B[1] & A[1]) | (B[2] & ~B[0] & A[1] & A[0]);
	assign D = (~B[2] & A[2]) | (~B[2] & B[0] & ~A[1] & ~A[0]) | (~B[2] & B[1] & ~A[1]) | (~B[2] & B[1] & B[0] & ~A[0]) | (B[0] & A[2] & ~A[1] & ~A[0]) | (B[1] & A[2] & ~A[1]) | (B[1] & B[0] & A[2] & ~A[0]);
endmodule
